module shift_left_4 (input [23:0] a, output [23:0] b);
  assign b = a << 4;
endmodule