module _1x8uExt (input in, output [7:0] out);
  assign out = {7'b0, in};
endmodule